LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY RECLAMA IS
	PORT( BUTON_IN: IN STD_LOGIC_VECTOR(2 DOWNTO 0);	
			WE: IN STD_LOGIC;
			ANIMATIE: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			CLK: IN STD_LOGIC;
			RESET: IN STD_LOGIC;
			AN: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			SEG: OUT STD_LOGIC_VECTOR(0 TO 7));
END ENTITY;

ARCHITECTURE ARCH_RECLAMA OF RECLAMA IS	  

SIGNAL BUTON_OUT: STD_LOGIC_VECTOR(2 DOWNTO 0); --BUTOANELE DUPA DEBOUNCE
SIGNAL T: STD_LOGIC; --NOUL CLOCK CU FRECVENTA DE 1 SECUNDA
SIGNAL S: STD_LOGIC; --CLOCK DIVIZAT PENTRU REGISTRU
SIGNAL TEMPO: STD_LOGIC_VECTOR(1 DOWNTO 0);	 --PENTRU SCHIMBARE ANODURILOR
SIGNAL Y: INTEGER RANGE 0 TO 3:=3; --PENTRU ALEGEREA LITERELOR
SIGNAL CONT: INTEGER RANGE 0 TO 4:=0; --PENTRU ALEGEREA LITERELOR
SIGNAL I: INTEGER RANGE 0 TO 4:=0; --PENTRU DEPLASARE
SIGNAL DATA1, DATA2, DATA3, DATA4 : STD_LOGIC_VECTOR(0 TO 7):="11111111"; --PENTRU DEPLASARE 
SIGNAL C1, C2, C3, C4 : STD_LOGIC_VECTOR(0 TO 7):="11111111"; --PENTRU PWM
SIGNAL D1, D2, D3, D4 : STD_LOGIC_VECTOR(0 TO 7):="11111111"; --PENTRU AFISARE LITERA CU LITERA
SIGNAL I1: INTEGER RANGE 0 TO 3:=0; --PENTRU AFISARE LITERA CU LITERA
SIGNAL COUNTER1: INTEGER RANGE 0 TO 2300; --PENTRU PWM
SIGNAL COUNTER2: INTEGER RANGE 0 TO 10500; --PENTRU PWM
SIGNAL VALOARE: INTEGER RANGE 0 TO 2300;	--PENTRU PWM
SIGNAL T1: STD_LOGIC; --PENTRU PWM
SIGNAL OK: STD_LOGIC; -- PENTRU PWM
TYPE MEMORIE1 IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE MEMORIE2 IS ARRAY (3 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

COMPONENT DIVIZOR1 IS 
PORT ( CLK : IN  STD_LOGIC;
       CLK_OUT : OUT STD_LOGIC);
END COMPONENT;

COMPONENT DIVIZOR2 IS 
PORT ( CLK : IN  STD_LOGIC;
       CLK_OUT : OUT STD_LOGIC);
END COMPONENT;

COMPONENT DEBOUNCE IS
PORT (CLK: IN STD_LOGIC;
		BUTON_IN : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		BUTON_OUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END COMPONENT;

COMPONENT DIVIZORAN IS 
PORT (CLK : IN STD_LOGIC;
		TEMPO: OUT STD_LOGIC_VECTOR(1 DOWNTO 0));
END COMPONENT;

--MEMORIA DE SIMBOLURI
CONSTANT SIMBOL: MEMORIE1:=(
0=> "00000011", --0
1=> "10011111", --1	
2=> "00100101", --2
3=> "00001101",	--3
4=> "10011001",	--4
5=> "01001001",	--5
6=> "01000001",	--6
7=> "00011111",	--7
8=> "00000001",	--8
9=> "00001001",	--9
10=> "00010001",--A
11=> "11000001",--b
12=> "01100011",--C
13=> "10000101",--d
14=> "01100001",--E
15=> "01110001", --F
16=> "01000011", --G
17=> "10010001", --H
18=> "11110011", --I
19=> "10000111", --J
20=> "01010001", --k
21=> "11100011", --L
22=> "11010101", --n
23=> "11000101", --o
24=> "00110001", --P
25=> "00011001", --q
26=> "11110101", --r
27=> "01001001", --S
28=> "11100001", --t
29=> "10000011", --U
30=> "10001001", --y
31=> "11111111"); --spatiu

--INITIALIZARE MEMORIE CUVANT
SIGNAL CUVINTE: MEMORIE2:=(
0=> SIMBOL(31),
1=> SIMBOL(31),	
2=> SIMBOL(31),
3=> SIMBOL(31));

BEGIN

--DEBOUNCE BUTOANE	
DEBOUNCEBUTOANE: DEBOUNCE PORT MAP (CLK, BUTON_IN, BUTON_OUT); 

--DIVIZAREA DE FRECVENTA PENTRU CLIPIRE
DIVIZOR1SEC: DIVIZOR1 PORT MAP (CLK,T);

--DIVIZOR PENTRU SCHIMBARE ANODURILOR
DIVIZORANODURI: DIVIZORAN PORT MAP (CLK, TEMPO);

--DIVIZOR PENTRU DEPLASARE
DIVIZORDEPLASARE: DIVIZOR2 PORT MAP (CLK,S);

--AFISAREA EFECTIVA
PROCESS(T, TEMPO, ANIMATIE, BUTON_OUT)
VARIABLE X: INTEGER RANGE 0 TO 31:=0;
BEGIN
--ALEGEREA LITERELOR DIN CUVANT
IF RESET='0' THEN
IF WE='1' THEN
			IF CONT=0 THEN
				AN<="1110";
				SEG<=SIMBOL(X);
			ELSIF CONT=1 THEN 
				IF TEMPO="00" OR TEMPO="10" THEN AN<="1110"; SEG<=SIMBOL(X);
				ELSE AN<="1101"; SEG<=CUVINTE(3);
				END IF;
			ELSIF CONT=2 THEN
				IF TEMPO="00" OR TEMPO="10" THEN AN<="1110"; SEG<=SIMBOL(X);
				ELSIF TEMPO="01" THEN  AN<="1101"; SEG<=CUVINTE(2);
				ELSE AN<="1011"; SEG<=CUVINTE(3);
				END IF;
			ELSIF CONT=3 THEN 
				IF TEMPO="00" THEN
					AN<="1110"; SEG<=SIMBOL(X);
				ELSIF TEMPO="01" THEN  AN<="1101"; SEG<=CUVINTE(1);
				ELSIF TEMPO="10" THEN AN<="1011"; SEG<=CUVINTE(2);
				ELSE AN<="0111"; SEG<=CUVINTE(3);
				END IF;
			ELSIF CONT=4 THEN
				IF TEMPO="00" THEN AN<="1110"; SEG<=CUVINTE(0);
				ELSIF TEMPO="01" THEN  AN<="1101"; SEG<=CUVINTE(1);
				ELSIF TEMPO="10" THEN AN<="1011"; SEG<=CUVINTE(2);
				ELSE AN<="0111"; SEG<=CUVINTE(3);
				END IF;
			END IF;
		
	IF RISING_EDGE(BUTON_OUT(1)) THEN X:=X+1;
	END IF;
	
	IF RISING_EDGE(BUTON_OUT(0)) THEN 
				IF CONT<4  THEN 
					CONT<=CONT+1;
					CUVINTE(Y)<=SIMBOL(X);
					Y<=Y-1;
				END IF;
	END IF;

ELSE 
--AFISAREA CUVANTULUI ALES
	IF ANIMATIE="000" OR ANIMATIE="101" OR ANIMATIE="110" OR ANIMATIE="111" THEN --AFISARE CONTINUA
		 CASE TEMPO IS
						WHEN "00" => AN<="1110"; SEG<=CUVINTE(0);
						WHEN "01" => AN<="1101"; SEG<=CUVINTE(1);
						WHEN "10" => AN<="1011"; SEG<=CUVINTE(2);
						WHEN "11" => AN<="0111"; SEG<=CUVINTE(3); 	
						WHEN OTHERS => AN<="1111"; SEG<=SIMBOL(14);
		END CASE;

	ELSIF ANIMATIE="001" THEN --CLIPIRE
		IF T='1' THEN
			CASE TEMPO IS
						WHEN "00" => AN<="1110"; SEG<=CUVINTE(0);
						WHEN "01" => AN<="1101"; SEG<=CUVINTE(1);
						WHEN "10" => AN<="1011"; SEG<=CUVINTE(2);
						WHEN "11" => AN<="0111"; SEG<=CUVINTE(3); 
						WHEN OTHERS => AN<="1111"; SEG<=SIMBOL(14);
			END CASE;
		ELSE AN<="1111";
		END IF;
	ELSIF ANIMATIE="010" THEN --DEPLASARE DREAPTA -> STANGA
		IF RISING_EDGE(S) THEN 
		--DEPLASARE (SE FACE CONCURENT);	
			IF I=4 THEN 
				DATA1<="11111111";
				DATA2<=DATA1;
				DATA3<=DATA2;
				DATA4<=DATA3;
				I<=0;
			ELSE 
				DATA1<=CUVINTE(3-I);
				DATA2<=DATA1;
				DATA3<=DATA2;
				DATA4<=DATA3;
				I<=I+1;
			END IF;
		END IF;
	
			CASE TEMPO IS
						WHEN "00" => AN<="1110"; SEG<=DATA1;
						WHEN "01" => AN<="1101"; SEG<=DATA2;
						WHEN "10" => AN<="1011"; SEG<=DATA3;
						WHEN "11" => AN<="0111"; SEG<=DATA4; 
						WHEN OTHERS => AN<="1111"; SEG<=SIMBOL(14);
			END CASE;	
	ELSIF ANIMATIE="011" THEN --INTENSITATE VARIABILA (PWM)
				
IF RISING_EDGE(CLK) THEN
	IF COUNTER1=2299 THEN --NUMARA CAT SA FIE APRINS 
	COUNTER1<=0;
	ELSE COUNTER1<=COUNTER1+1;
	END IF;
	
	IF COUNTER1<=VALOARE THEN 
	C1<=CUVINTE(0);
	C2<=CUVINTE(1);
	C3<=CUVINTE(2);
	C4<=CUVINTE(3);
	ELSE 
	C1<="11111111";
	C2<="11111111";
	C3<="11111111";
	C4<="11111111";
	END IF;
	
	IF COUNTER2=10499 THEN --DIVIZEAZA CLOCK-UL PENTRU A DETERMINA MODIFICAREA VALORII CURENTE
		COUNTER2<=0;
		T1<=NOT T1;
	ELSE COUNTER2<=COUNTER2+1;
	END IF;
	
END IF;

IF RISING_EDGE(T1) THEN 
	IF OK='0' AND VALOARE<2299 THEN VALOARE<=VALOARE+1;
	ELSIF OK='0' AND VALOARE>=2299 THEN OK<='1'; VALOARE<=VALOARE-1;
	ELSIF OK='1' AND VALOARE>0 THEN VALOARE<=VALOARE-1;
	ELSIF OK='1' AND VALOARE=0 THEN OK<='0'; VALOARE<=VALOARE+1;
	END IF;
END IF;

			CASE TEMPO IS
						WHEN "00" => AN<="1110"; SEG<=C1;
						WHEN "01" => AN<="1101"; SEG<=C2;
						WHEN "10" => AN<="1011"; SEG<=C3;
						WHEN "11" => AN<="0111"; SEG<=C4; 
						WHEN OTHERS => AN<="1111"; SEG<=SIMBOL(14);
			END CASE;	

ELSIF ANIMATIE="100" THEN --AFISARE LITERA CU LITERA 

IF RISING_EDGE(S) THEN 
		--DEPLASARE (SE FACE CONCURENT);	
		IF I1=0 THEN 
			D1<=CUVINTE(3);
			D2<="11111101";
			D3<="11111101";
			D4<="11111101";
		ELSIF I1=1 THEN 
			D1<="11111101";
			D2<=CUVINTE(2);
			D3<="11111101";
			D4<="11111101";
		ELSIF I1=2 THEN 
			D1<="11111101";
			D2<="11111101";
			D3<=CUVINTE(1);
			D4<="11111101";
		ELSIF I1=3 THEN 
			D1<="11111101";
			D2<="11111101";
			D3<="11111101";
			D4<=CUVINTE(0);
		END IF;
		
		IF I1<3 THEN I1<=I1+1;
		ELSE I1<=0;
		END IF;
		
	END IF;
		CASE TEMPO IS
						WHEN "00" => AN<="1110"; SEG<=D4;
						WHEN "01" => AN<="1101"; SEG<=D3;
						WHEN "10" => AN<="1011"; SEG<=D2;
						WHEN "11" => AN<="0111"; SEG<=D1; 
						WHEN OTHERS => AN<="1111"; SEG<=SIMBOL(14);
			END CASE;
END IF; --IF DE LA ANIMATIE
END IF; --IF DE LA WE
ELSE 
	Y<=3;
	X:=0;
	CONT<=0;
	I<=0;
	I1<=0;
	DATA1<="11111111";
	DATA2<="11111111";
	DATA3<="11111111";
	DATA4<="11111111";
	C1<="11111111";
	C2<="11111111";
	C3<="11111111";
	C4<="11111111";
	D1<="11111111";
	D2<="11111111";
	D3<="11111111";
	D4<="11111111";
	SEG<="11111111";
	AN<="1111";
	CUVINTE(0)<="11111111";
	CUVINTE(1)<="11111111";
	CUVINTE(2)<="11111111";
	CUVINTE(3)<="11111111";
END IF; --IF DE LA RESET		
END PROCESS;
END ARCHITECTURE;