LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DIVIZOR1 IS 
	PORT (CLK: IN STD_LOGIC;
			CLK_OUT: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE ARCH_DIVIZOR1 OF DIVIZOR1 IS
SIGNAL COUNTER_DIV: INTEGER RANGE 0 TO 25000000:=0;
SIGNAL T: STD_LOGIC;
BEGIN
PROCESS(CLK)
BEGIN
	IF RISING_EDGE(CLK) THEN 
		IF COUNTER_DIV=24999999 THEN 
			COUNTER_DIV<=0;
			T<=NOT T;
		ELSE COUNTER_DIV<=COUNTER_DIV+1;
		END IF;
	END IF;
END PROCESS;
CLK_OUT<=T;
END ARCHITECTURE;