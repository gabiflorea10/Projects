LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DIVIZOR2 IS 
	PORT (CLK: IN STD_LOGIC;
			CLK_OUT: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE ARCH_DIVIZOR2 OF DIVIZOR2 IS
SIGNAL COUNTER_DIV: INTEGER RANGE 0 TO 18000000:=0;
SIGNAL S: STD_LOGIC;
BEGIN
PROCESS(CLK)
BEGIN
	IF RISING_EDGE(CLK) THEN 
		IF COUNTER_DIV=17999999 THEN 
			COUNTER_DIV<=0;
			S<=NOT S;
		ELSE COUNTER_DIV<=COUNTER_DIV+1;
		END IF;
	END IF;
END PROCESS;
CLK_OUT<=S;
END ARCHITECTURE;