LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEBOUNCE IS
	PORT( CLK: IN STD_LOGIC;
			BUTON_IN: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			BUTON_OUT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END ENTITY;

ARCHITECTURE ARCH_DEBOUNCE OF DEBOUNCE IS
SIGNAL COUNTER: INTEGER RANGE 0 TO 500000:=0;
SIGNAL D1,D2,D3: STD_LOGIC_VECTOR (2 DOWNTO 0);
BEGIN
PROCESS(CLK)
BEGIN
	IF RISING_EDGE(CLK) THEN
		IF COUNTER=499999 THEN 
			COUNTER<=0;
			D1<=BUTON_IN;
			D2<=D1;
			D3<=D2;
		ELSE COUNTER<=COUNTER+1;
		END IF;
	END IF;
END PROCESS;
BUTON_OUT<=D1 AND D2 AND D3;
END ARCHITECTURE;